module adder (
    input [19:0] a,
    input [19:0] b,
    output [19:0] sum
);
    assign sum = a + b;
endmodule

